`default_nettype none

module spi_peripheral(
    input wire COPI,
    input wire nCS,
    input wire SCLK,

);


endmodule